module Rcon(
	input wire [3:0] j,
	output wire [31:0] Rcon_j
);
	assign Rcon_j = (j == 4'b0001) ? 32'h01000000 :
						 (j == 4'b0010) ? 32'h02000000 :
						 (j == 4'b0011) ? 32'h04000000 :
						 (j == 4'b0100) ? 32'h08000000 :
						 (j == 4'b0101) ? 32'h10000000 :
						 (j == 4'b0110) ? 32'h20000000 :
						 (j == 4'b0111) ? 32'h40000000 :
						 (j == 4'b1000) ? 32'h80000000 :
						 (j == 4'b1001) ? 32'h1b000000 :
						 (j == 4'b1010) ? 32'h36000000 :
						  32'b0; // Default case
endmodule
